module libretrov

pub const (
	retro_api_version = 1
	retro_num_core_options_values_max = 128
)